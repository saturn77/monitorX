// NiosBase.v

// Generated using ACDS version 20.1 720

`timescale 1 ps / 1 ps
module NiosBase (
		input  wire        clk_clk,           //        clk.clk
		input  wire        coe_done,          //        coe.done
		input  wire [7:0]  coe_data,          //           .data
		input  wire [15:0] i_reg16_0_export,  //  i_reg16_0.export
		input  wire [15:0] i_reg16_1_export,  //  i_reg16_1.export
		input  wire [15:0] i_reg16_2_export,  //  i_reg16_2.export
		input  wire [15:0] i_reg16_3_export,  //  i_reg16_3.export
		input  wire [15:0] i_reg16_4_export,  //  i_reg16_4.export
		input  wire [15:0] i_reg16_5_export,  //  i_reg16_5.export
		input  wire [15:0] i_reg16_6_export,  //  i_reg16_6.export
		input  wire [31:0] i_reg32_0_export,  //  i_reg32_0.export
		input  wire [31:0] i_reg32_1_export,  //  i_reg32_1.export
		input  wire [31:0] i_reg32_2_export,  //  i_reg32_2.export
		input  wire [31:0] i_reg32_3_export,  //  i_reg32_3.export
		input  wire [31:0] i_reg32_4_export,  //  i_reg32_4.export
		input  wire [31:0] i_reg32_5_export,  //  i_reg32_5.export
		input  wire [31:0] i_reg32_6_export,  //  i_reg32_6.export
		input  wire [31:0] i_reg32_7_export,  //  i_reg32_7.export
		output wire [31:0] o_reg32_0_export,  //  o_reg32_0.export
		output wire [31:0] o_reg32_1_export,  //  o_reg32_1.export
		output wire [31:0] o_reg32_10_export, // o_reg32_10.export
		output wire [31:0] o_reg32_11_export, // o_reg32_11.export
		output wire [31:0] o_reg32_12_export, // o_reg32_12.export
		output wire [31:0] o_reg32_13_export, // o_reg32_13.export
		output wire [31:0] o_reg32_2_export,  //  o_reg32_2.export
		output wire [31:0] o_reg32_3_export,  //  o_reg32_3.export
		output wire [31:0] o_reg32_4_export,  //  o_reg32_4.export
		output wire [31:0] o_reg32_5_export,  //  o_reg32_5.export
		output wire [31:0] o_reg32_6_export,  //  o_reg32_6.export
		output wire [31:0] o_reg32_7_export,  //  o_reg32_7.export
		output wire [31:0] o_reg32_8_export,  //  o_reg32_8.export
		output wire [31:0] o_reg32_9_export,  //  o_reg32_9.export
		input  wire        reset_reset_n,     //      reset.reset_n
		input  wire        uart_rxd,          //       uart.rxd
		output wire        uart_txd           //           .txd
	);

	wire  [31:0] nios2_gen2_0_data_master_readdata;                          // mm_interconnect_0:nios2_gen2_0_data_master_readdata -> nios2_gen2_0:d_readdata
	wire         nios2_gen2_0_data_master_waitrequest;                       // mm_interconnect_0:nios2_gen2_0_data_master_waitrequest -> nios2_gen2_0:d_waitrequest
	wire         nios2_gen2_0_data_master_debugaccess;                       // nios2_gen2_0:debug_mem_slave_debugaccess_to_roms -> mm_interconnect_0:nios2_gen2_0_data_master_debugaccess
	wire  [18:0] nios2_gen2_0_data_master_address;                           // nios2_gen2_0:d_address -> mm_interconnect_0:nios2_gen2_0_data_master_address
	wire   [3:0] nios2_gen2_0_data_master_byteenable;                        // nios2_gen2_0:d_byteenable -> mm_interconnect_0:nios2_gen2_0_data_master_byteenable
	wire         nios2_gen2_0_data_master_read;                              // nios2_gen2_0:d_read -> mm_interconnect_0:nios2_gen2_0_data_master_read
	wire         nios2_gen2_0_data_master_write;                             // nios2_gen2_0:d_write -> mm_interconnect_0:nios2_gen2_0_data_master_write
	wire  [31:0] nios2_gen2_0_data_master_writedata;                         // nios2_gen2_0:d_writedata -> mm_interconnect_0:nios2_gen2_0_data_master_writedata
	wire  [31:0] nios2_gen2_0_instruction_master_readdata;                   // mm_interconnect_0:nios2_gen2_0_instruction_master_readdata -> nios2_gen2_0:i_readdata
	wire         nios2_gen2_0_instruction_master_waitrequest;                // mm_interconnect_0:nios2_gen2_0_instruction_master_waitrequest -> nios2_gen2_0:i_waitrequest
	wire  [18:0] nios2_gen2_0_instruction_master_address;                    // nios2_gen2_0:i_address -> mm_interconnect_0:nios2_gen2_0_instruction_master_address
	wire         nios2_gen2_0_instruction_master_read;                       // nios2_gen2_0:i_read -> mm_interconnect_0:nios2_gen2_0_instruction_master_read
	wire  [31:0] mm_interconnect_0_dma_rx_0_av_mm_readdata;                  // dma_rx_0:av_mm_readdata -> mm_interconnect_0:dma_rx_0_av_mm_readdata
	wire         mm_interconnect_0_dma_rx_0_av_mm_waitrequest;               // dma_rx_0:av_mm_waitrequest -> mm_interconnect_0:dma_rx_0_av_mm_waitrequest
	wire   [4:0] mm_interconnect_0_dma_rx_0_av_mm_address;                   // mm_interconnect_0:dma_rx_0_av_mm_address -> dma_rx_0:av_mm_addr
	wire         mm_interconnect_0_dma_rx_0_av_mm_read;                      // mm_interconnect_0:dma_rx_0_av_mm_read -> dma_rx_0:av_mm_read
	wire         mm_interconnect_0_dma_rx_0_av_mm_write;                     // mm_interconnect_0:dma_rx_0_av_mm_write -> dma_rx_0:av_mm_write
	wire  [31:0] mm_interconnect_0_dma_rx_0_av_mm_writedata;                 // mm_interconnect_0:dma_rx_0_av_mm_writedata -> dma_rx_0:av_mm_writedata
	wire  [31:0] mm_interconnect_0_nios2_gen2_0_debug_mem_slave_readdata;    // nios2_gen2_0:debug_mem_slave_readdata -> mm_interconnect_0:nios2_gen2_0_debug_mem_slave_readdata
	wire         mm_interconnect_0_nios2_gen2_0_debug_mem_slave_waitrequest; // nios2_gen2_0:debug_mem_slave_waitrequest -> mm_interconnect_0:nios2_gen2_0_debug_mem_slave_waitrequest
	wire         mm_interconnect_0_nios2_gen2_0_debug_mem_slave_debugaccess; // mm_interconnect_0:nios2_gen2_0_debug_mem_slave_debugaccess -> nios2_gen2_0:debug_mem_slave_debugaccess
	wire   [8:0] mm_interconnect_0_nios2_gen2_0_debug_mem_slave_address;     // mm_interconnect_0:nios2_gen2_0_debug_mem_slave_address -> nios2_gen2_0:debug_mem_slave_address
	wire         mm_interconnect_0_nios2_gen2_0_debug_mem_slave_read;        // mm_interconnect_0:nios2_gen2_0_debug_mem_slave_read -> nios2_gen2_0:debug_mem_slave_read
	wire   [3:0] mm_interconnect_0_nios2_gen2_0_debug_mem_slave_byteenable;  // mm_interconnect_0:nios2_gen2_0_debug_mem_slave_byteenable -> nios2_gen2_0:debug_mem_slave_byteenable
	wire         mm_interconnect_0_nios2_gen2_0_debug_mem_slave_write;       // mm_interconnect_0:nios2_gen2_0_debug_mem_slave_write -> nios2_gen2_0:debug_mem_slave_write
	wire  [31:0] mm_interconnect_0_nios2_gen2_0_debug_mem_slave_writedata;   // mm_interconnect_0:nios2_gen2_0_debug_mem_slave_writedata -> nios2_gen2_0:debug_mem_slave_writedata
	wire         mm_interconnect_0_onchip_memory2_0_s1_chipselect;           // mm_interconnect_0:onchip_memory2_0_s1_chipselect -> onchip_memory2_0:chipselect
	wire  [31:0] mm_interconnect_0_onchip_memory2_0_s1_readdata;             // onchip_memory2_0:readdata -> mm_interconnect_0:onchip_memory2_0_s1_readdata
	wire  [14:0] mm_interconnect_0_onchip_memory2_0_s1_address;              // mm_interconnect_0:onchip_memory2_0_s1_address -> onchip_memory2_0:address
	wire   [3:0] mm_interconnect_0_onchip_memory2_0_s1_byteenable;           // mm_interconnect_0:onchip_memory2_0_s1_byteenable -> onchip_memory2_0:byteenable
	wire         mm_interconnect_0_onchip_memory2_0_s1_write;                // mm_interconnect_0:onchip_memory2_0_s1_write -> onchip_memory2_0:write
	wire  [31:0] mm_interconnect_0_onchip_memory2_0_s1_writedata;            // mm_interconnect_0:onchip_memory2_0_s1_writedata -> onchip_memory2_0:writedata
	wire         mm_interconnect_0_onchip_memory2_0_s1_clken;                // mm_interconnect_0:onchip_memory2_0_s1_clken -> onchip_memory2_0:clken
	wire         mm_interconnect_0_timer_0_s1_chipselect;                    // mm_interconnect_0:timer_0_s1_chipselect -> timer_0:chipselect
	wire  [15:0] mm_interconnect_0_timer_0_s1_readdata;                      // timer_0:readdata -> mm_interconnect_0:timer_0_s1_readdata
	wire   [2:0] mm_interconnect_0_timer_0_s1_address;                       // mm_interconnect_0:timer_0_s1_address -> timer_0:address
	wire         mm_interconnect_0_timer_0_s1_write;                         // mm_interconnect_0:timer_0_s1_write -> timer_0:write_n
	wire  [15:0] mm_interconnect_0_timer_0_s1_writedata;                     // mm_interconnect_0:timer_0_s1_writedata -> timer_0:writedata
	wire         mm_interconnect_0_timer_1_s1_chipselect;                    // mm_interconnect_0:timer_1_s1_chipselect -> timer_1:chipselect
	wire  [15:0] mm_interconnect_0_timer_1_s1_readdata;                      // timer_1:readdata -> mm_interconnect_0:timer_1_s1_readdata
	wire   [2:0] mm_interconnect_0_timer_1_s1_address;                       // mm_interconnect_0:timer_1_s1_address -> timer_1:address
	wire         mm_interconnect_0_timer_1_s1_write;                         // mm_interconnect_0:timer_1_s1_write -> timer_1:write_n
	wire  [15:0] mm_interconnect_0_timer_1_s1_writedata;                     // mm_interconnect_0:timer_1_s1_writedata -> timer_1:writedata
	wire         mm_interconnect_0_i_reg32_0_s1_chipselect;                  // mm_interconnect_0:i_reg32_0_s1_chipselect -> i_reg32_0:chipselect
	wire  [31:0] mm_interconnect_0_i_reg32_0_s1_readdata;                    // i_reg32_0:readdata -> mm_interconnect_0:i_reg32_0_s1_readdata
	wire   [1:0] mm_interconnect_0_i_reg32_0_s1_address;                     // mm_interconnect_0:i_reg32_0_s1_address -> i_reg32_0:address
	wire         mm_interconnect_0_i_reg32_0_s1_write;                       // mm_interconnect_0:i_reg32_0_s1_write -> i_reg32_0:write_n
	wire  [31:0] mm_interconnect_0_i_reg32_0_s1_writedata;                   // mm_interconnect_0:i_reg32_0_s1_writedata -> i_reg32_0:writedata
	wire  [31:0] mm_interconnect_0_i_reg32_1_s1_readdata;                    // i_reg32_1:readdata -> mm_interconnect_0:i_reg32_1_s1_readdata
	wire   [1:0] mm_interconnect_0_i_reg32_1_s1_address;                     // mm_interconnect_0:i_reg32_1_s1_address -> i_reg32_1:address
	wire  [31:0] mm_interconnect_0_i_reg16_0_s1_readdata;                    // i_reg16_0:readdata -> mm_interconnect_0:i_reg16_0_s1_readdata
	wire   [1:0] mm_interconnect_0_i_reg16_0_s1_address;                     // mm_interconnect_0:i_reg16_0_s1_address -> i_reg16_0:address
	wire  [31:0] mm_interconnect_0_i_reg16_1_s1_readdata;                    // i_reg16_1:readdata -> mm_interconnect_0:i_reg16_1_s1_readdata
	wire   [1:0] mm_interconnect_0_i_reg16_1_s1_address;                     // mm_interconnect_0:i_reg16_1_s1_address -> i_reg16_1:address
	wire  [31:0] mm_interconnect_0_i_reg16_2_s1_readdata;                    // i_reg16_2:readdata -> mm_interconnect_0:i_reg16_2_s1_readdata
	wire   [1:0] mm_interconnect_0_i_reg16_2_s1_address;                     // mm_interconnect_0:i_reg16_2_s1_address -> i_reg16_2:address
	wire  [31:0] mm_interconnect_0_i_reg16_3_s1_readdata;                    // i_reg16_3:readdata -> mm_interconnect_0:i_reg16_3_s1_readdata
	wire   [1:0] mm_interconnect_0_i_reg16_3_s1_address;                     // mm_interconnect_0:i_reg16_3_s1_address -> i_reg16_3:address
	wire  [31:0] mm_interconnect_0_i_reg16_4_s1_readdata;                    // i_reg16_4:readdata -> mm_interconnect_0:i_reg16_4_s1_readdata
	wire   [1:0] mm_interconnect_0_i_reg16_4_s1_address;                     // mm_interconnect_0:i_reg16_4_s1_address -> i_reg16_4:address
	wire  [31:0] mm_interconnect_0_i_reg16_5_s1_readdata;                    // i_reg16_5:readdata -> mm_interconnect_0:i_reg16_5_s1_readdata
	wire   [1:0] mm_interconnect_0_i_reg16_5_s1_address;                     // mm_interconnect_0:i_reg16_5_s1_address -> i_reg16_5:address
	wire  [31:0] mm_interconnect_0_i_reg16_6_s1_readdata;                    // i_reg16_6:readdata -> mm_interconnect_0:i_reg16_6_s1_readdata
	wire   [1:0] mm_interconnect_0_i_reg16_6_s1_address;                     // mm_interconnect_0:i_reg16_6_s1_address -> i_reg16_6:address
	wire         mm_interconnect_0_uart_0_s1_chipselect;                     // mm_interconnect_0:uart_0_s1_chipselect -> uart_0:chipselect
	wire  [15:0] mm_interconnect_0_uart_0_s1_readdata;                       // uart_0:readdata -> mm_interconnect_0:uart_0_s1_readdata
	wire   [2:0] mm_interconnect_0_uart_0_s1_address;                        // mm_interconnect_0:uart_0_s1_address -> uart_0:address
	wire         mm_interconnect_0_uart_0_s1_read;                           // mm_interconnect_0:uart_0_s1_read -> uart_0:read_n
	wire         mm_interconnect_0_uart_0_s1_begintransfer;                  // mm_interconnect_0:uart_0_s1_begintransfer -> uart_0:begintransfer
	wire         mm_interconnect_0_uart_0_s1_write;                          // mm_interconnect_0:uart_0_s1_write -> uart_0:write_n
	wire  [15:0] mm_interconnect_0_uart_0_s1_writedata;                      // mm_interconnect_0:uart_0_s1_writedata -> uart_0:writedata
	wire         mm_interconnect_0_o_reg32_0_s1_chipselect;                  // mm_interconnect_0:o_reg32_0_s1_chipselect -> o_reg32_0:chipselect
	wire  [31:0] mm_interconnect_0_o_reg32_0_s1_readdata;                    // o_reg32_0:readdata -> mm_interconnect_0:o_reg32_0_s1_readdata
	wire   [1:0] mm_interconnect_0_o_reg32_0_s1_address;                     // mm_interconnect_0:o_reg32_0_s1_address -> o_reg32_0:address
	wire         mm_interconnect_0_o_reg32_0_s1_write;                       // mm_interconnect_0:o_reg32_0_s1_write -> o_reg32_0:write_n
	wire  [31:0] mm_interconnect_0_o_reg32_0_s1_writedata;                   // mm_interconnect_0:o_reg32_0_s1_writedata -> o_reg32_0:writedata
	wire         mm_interconnect_0_o_reg32_1_s1_chipselect;                  // mm_interconnect_0:o_reg32_1_s1_chipselect -> o_reg32_1:chipselect
	wire  [31:0] mm_interconnect_0_o_reg32_1_s1_readdata;                    // o_reg32_1:readdata -> mm_interconnect_0:o_reg32_1_s1_readdata
	wire   [1:0] mm_interconnect_0_o_reg32_1_s1_address;                     // mm_interconnect_0:o_reg32_1_s1_address -> o_reg32_1:address
	wire         mm_interconnect_0_o_reg32_1_s1_write;                       // mm_interconnect_0:o_reg32_1_s1_write -> o_reg32_1:write_n
	wire  [31:0] mm_interconnect_0_o_reg32_1_s1_writedata;                   // mm_interconnect_0:o_reg32_1_s1_writedata -> o_reg32_1:writedata
	wire         mm_interconnect_0_o_reg32_2_s1_chipselect;                  // mm_interconnect_0:o_reg32_2_s1_chipselect -> o_reg32_2:chipselect
	wire  [31:0] mm_interconnect_0_o_reg32_2_s1_readdata;                    // o_reg32_2:readdata -> mm_interconnect_0:o_reg32_2_s1_readdata
	wire   [1:0] mm_interconnect_0_o_reg32_2_s1_address;                     // mm_interconnect_0:o_reg32_2_s1_address -> o_reg32_2:address
	wire         mm_interconnect_0_o_reg32_2_s1_write;                       // mm_interconnect_0:o_reg32_2_s1_write -> o_reg32_2:write_n
	wire  [31:0] mm_interconnect_0_o_reg32_2_s1_writedata;                   // mm_interconnect_0:o_reg32_2_s1_writedata -> o_reg32_2:writedata
	wire         mm_interconnect_0_o_reg32_3_s1_chipselect;                  // mm_interconnect_0:o_reg32_3_s1_chipselect -> o_reg32_3:chipselect
	wire  [31:0] mm_interconnect_0_o_reg32_3_s1_readdata;                    // o_reg32_3:readdata -> mm_interconnect_0:o_reg32_3_s1_readdata
	wire   [1:0] mm_interconnect_0_o_reg32_3_s1_address;                     // mm_interconnect_0:o_reg32_3_s1_address -> o_reg32_3:address
	wire         mm_interconnect_0_o_reg32_3_s1_write;                       // mm_interconnect_0:o_reg32_3_s1_write -> o_reg32_3:write_n
	wire  [31:0] mm_interconnect_0_o_reg32_3_s1_writedata;                   // mm_interconnect_0:o_reg32_3_s1_writedata -> o_reg32_3:writedata
	wire         mm_interconnect_0_o_reg32_4_s1_chipselect;                  // mm_interconnect_0:o_reg32_4_s1_chipselect -> o_reg32_4:chipselect
	wire  [31:0] mm_interconnect_0_o_reg32_4_s1_readdata;                    // o_reg32_4:readdata -> mm_interconnect_0:o_reg32_4_s1_readdata
	wire   [1:0] mm_interconnect_0_o_reg32_4_s1_address;                     // mm_interconnect_0:o_reg32_4_s1_address -> o_reg32_4:address
	wire         mm_interconnect_0_o_reg32_4_s1_write;                       // mm_interconnect_0:o_reg32_4_s1_write -> o_reg32_4:write_n
	wire  [31:0] mm_interconnect_0_o_reg32_4_s1_writedata;                   // mm_interconnect_0:o_reg32_4_s1_writedata -> o_reg32_4:writedata
	wire         mm_interconnect_0_o_reg32_5_s1_chipselect;                  // mm_interconnect_0:o_reg32_5_s1_chipselect -> o_reg32_5:chipselect
	wire  [31:0] mm_interconnect_0_o_reg32_5_s1_readdata;                    // o_reg32_5:readdata -> mm_interconnect_0:o_reg32_5_s1_readdata
	wire   [1:0] mm_interconnect_0_o_reg32_5_s1_address;                     // mm_interconnect_0:o_reg32_5_s1_address -> o_reg32_5:address
	wire         mm_interconnect_0_o_reg32_5_s1_write;                       // mm_interconnect_0:o_reg32_5_s1_write -> o_reg32_5:write_n
	wire  [31:0] mm_interconnect_0_o_reg32_5_s1_writedata;                   // mm_interconnect_0:o_reg32_5_s1_writedata -> o_reg32_5:writedata
	wire         mm_interconnect_0_o_reg32_6_s1_chipselect;                  // mm_interconnect_0:o_reg32_6_s1_chipselect -> o_reg32_6:chipselect
	wire  [31:0] mm_interconnect_0_o_reg32_6_s1_readdata;                    // o_reg32_6:readdata -> mm_interconnect_0:o_reg32_6_s1_readdata
	wire   [1:0] mm_interconnect_0_o_reg32_6_s1_address;                     // mm_interconnect_0:o_reg32_6_s1_address -> o_reg32_6:address
	wire         mm_interconnect_0_o_reg32_6_s1_write;                       // mm_interconnect_0:o_reg32_6_s1_write -> o_reg32_6:write_n
	wire  [31:0] mm_interconnect_0_o_reg32_6_s1_writedata;                   // mm_interconnect_0:o_reg32_6_s1_writedata -> o_reg32_6:writedata
	wire         mm_interconnect_0_o_reg32_7_s1_chipselect;                  // mm_interconnect_0:o_reg32_7_s1_chipselect -> o_reg32_7:chipselect
	wire  [31:0] mm_interconnect_0_o_reg32_7_s1_readdata;                    // o_reg32_7:readdata -> mm_interconnect_0:o_reg32_7_s1_readdata
	wire   [1:0] mm_interconnect_0_o_reg32_7_s1_address;                     // mm_interconnect_0:o_reg32_7_s1_address -> o_reg32_7:address
	wire         mm_interconnect_0_o_reg32_7_s1_write;                       // mm_interconnect_0:o_reg32_7_s1_write -> o_reg32_7:write_n
	wire  [31:0] mm_interconnect_0_o_reg32_7_s1_writedata;                   // mm_interconnect_0:o_reg32_7_s1_writedata -> o_reg32_7:writedata
	wire         mm_interconnect_0_o_reg32_8_s1_chipselect;                  // mm_interconnect_0:o_reg32_8_s1_chipselect -> o_reg32_8:chipselect
	wire  [31:0] mm_interconnect_0_o_reg32_8_s1_readdata;                    // o_reg32_8:readdata -> mm_interconnect_0:o_reg32_8_s1_readdata
	wire   [1:0] mm_interconnect_0_o_reg32_8_s1_address;                     // mm_interconnect_0:o_reg32_8_s1_address -> o_reg32_8:address
	wire         mm_interconnect_0_o_reg32_8_s1_write;                       // mm_interconnect_0:o_reg32_8_s1_write -> o_reg32_8:write_n
	wire  [31:0] mm_interconnect_0_o_reg32_8_s1_writedata;                   // mm_interconnect_0:o_reg32_8_s1_writedata -> o_reg32_8:writedata
	wire         mm_interconnect_0_o_reg32_9_s1_chipselect;                  // mm_interconnect_0:o_reg32_9_s1_chipselect -> o_reg32_9:chipselect
	wire  [31:0] mm_interconnect_0_o_reg32_9_s1_readdata;                    // o_reg32_9:readdata -> mm_interconnect_0:o_reg32_9_s1_readdata
	wire   [1:0] mm_interconnect_0_o_reg32_9_s1_address;                     // mm_interconnect_0:o_reg32_9_s1_address -> o_reg32_9:address
	wire         mm_interconnect_0_o_reg32_9_s1_write;                       // mm_interconnect_0:o_reg32_9_s1_write -> o_reg32_9:write_n
	wire  [31:0] mm_interconnect_0_o_reg32_9_s1_writedata;                   // mm_interconnect_0:o_reg32_9_s1_writedata -> o_reg32_9:writedata
	wire         mm_interconnect_0_o_reg32_10_s1_chipselect;                 // mm_interconnect_0:o_reg32_10_s1_chipselect -> o_reg32_10:chipselect
	wire  [31:0] mm_interconnect_0_o_reg32_10_s1_readdata;                   // o_reg32_10:readdata -> mm_interconnect_0:o_reg32_10_s1_readdata
	wire   [1:0] mm_interconnect_0_o_reg32_10_s1_address;                    // mm_interconnect_0:o_reg32_10_s1_address -> o_reg32_10:address
	wire         mm_interconnect_0_o_reg32_10_s1_write;                      // mm_interconnect_0:o_reg32_10_s1_write -> o_reg32_10:write_n
	wire  [31:0] mm_interconnect_0_o_reg32_10_s1_writedata;                  // mm_interconnect_0:o_reg32_10_s1_writedata -> o_reg32_10:writedata
	wire         mm_interconnect_0_o_reg32_11_s1_chipselect;                 // mm_interconnect_0:o_reg32_11_s1_chipselect -> o_reg32_11:chipselect
	wire  [31:0] mm_interconnect_0_o_reg32_11_s1_readdata;                   // o_reg32_11:readdata -> mm_interconnect_0:o_reg32_11_s1_readdata
	wire   [1:0] mm_interconnect_0_o_reg32_11_s1_address;                    // mm_interconnect_0:o_reg32_11_s1_address -> o_reg32_11:address
	wire         mm_interconnect_0_o_reg32_11_s1_write;                      // mm_interconnect_0:o_reg32_11_s1_write -> o_reg32_11:write_n
	wire  [31:0] mm_interconnect_0_o_reg32_11_s1_writedata;                  // mm_interconnect_0:o_reg32_11_s1_writedata -> o_reg32_11:writedata
	wire  [31:0] mm_interconnect_0_i_reg32_2_s1_readdata;                    // i_reg32_2:readdata -> mm_interconnect_0:i_reg32_2_s1_readdata
	wire   [1:0] mm_interconnect_0_i_reg32_2_s1_address;                     // mm_interconnect_0:i_reg32_2_s1_address -> i_reg32_2:address
	wire  [31:0] mm_interconnect_0_i_reg32_3_s1_readdata;                    // i_reg32_3:readdata -> mm_interconnect_0:i_reg32_3_s1_readdata
	wire   [1:0] mm_interconnect_0_i_reg32_3_s1_address;                     // mm_interconnect_0:i_reg32_3_s1_address -> i_reg32_3:address
	wire  [31:0] mm_interconnect_0_i_reg32_4_s1_readdata;                    // i_reg32_4:readdata -> mm_interconnect_0:i_reg32_4_s1_readdata
	wire   [1:0] mm_interconnect_0_i_reg32_4_s1_address;                     // mm_interconnect_0:i_reg32_4_s1_address -> i_reg32_4:address
	wire  [31:0] mm_interconnect_0_i_reg32_5_s1_readdata;                    // i_reg32_5:readdata -> mm_interconnect_0:i_reg32_5_s1_readdata
	wire   [1:0] mm_interconnect_0_i_reg32_5_s1_address;                     // mm_interconnect_0:i_reg32_5_s1_address -> i_reg32_5:address
	wire  [31:0] mm_interconnect_0_i_reg32_6_s1_readdata;                    // i_reg32_6:readdata -> mm_interconnect_0:i_reg32_6_s1_readdata
	wire   [1:0] mm_interconnect_0_i_reg32_6_s1_address;                     // mm_interconnect_0:i_reg32_6_s1_address -> i_reg32_6:address
	wire  [31:0] mm_interconnect_0_i_reg32_7_s1_readdata;                    // i_reg32_7:readdata -> mm_interconnect_0:i_reg32_7_s1_readdata
	wire   [1:0] mm_interconnect_0_i_reg32_7_s1_address;                     // mm_interconnect_0:i_reg32_7_s1_address -> i_reg32_7:address
	wire         mm_interconnect_0_o_reg32_13_s1_chipselect;                 // mm_interconnect_0:o_reg32_13_s1_chipselect -> o_reg32_13:chipselect
	wire  [31:0] mm_interconnect_0_o_reg32_13_s1_readdata;                   // o_reg32_13:readdata -> mm_interconnect_0:o_reg32_13_s1_readdata
	wire   [1:0] mm_interconnect_0_o_reg32_13_s1_address;                    // mm_interconnect_0:o_reg32_13_s1_address -> o_reg32_13:address
	wire         mm_interconnect_0_o_reg32_13_s1_write;                      // mm_interconnect_0:o_reg32_13_s1_write -> o_reg32_13:write_n
	wire  [31:0] mm_interconnect_0_o_reg32_13_s1_writedata;                  // mm_interconnect_0:o_reg32_13_s1_writedata -> o_reg32_13:writedata
	wire         mm_interconnect_0_o_reg32_12_s1_chipselect;                 // mm_interconnect_0:o_reg32_12_s1_chipselect -> o_reg32_12:chipselect
	wire  [31:0] mm_interconnect_0_o_reg32_12_s1_readdata;                   // o_reg32_12:readdata -> mm_interconnect_0:o_reg32_12_s1_readdata
	wire   [1:0] mm_interconnect_0_o_reg32_12_s1_address;                    // mm_interconnect_0:o_reg32_12_s1_address -> o_reg32_12:address
	wire         mm_interconnect_0_o_reg32_12_s1_write;                      // mm_interconnect_0:o_reg32_12_s1_write -> o_reg32_12:write_n
	wire  [31:0] mm_interconnect_0_o_reg32_12_s1_writedata;                  // mm_interconnect_0:o_reg32_12_s1_writedata -> o_reg32_12:writedata
	wire         irq_mapper_receiver0_irq;                                   // timer_0:irq -> irq_mapper:receiver0_irq
	wire         irq_mapper_receiver1_irq;                                   // timer_1:irq -> irq_mapper:receiver1_irq
	wire         irq_mapper_receiver2_irq;                                   // i_reg32_0:irq -> irq_mapper:receiver2_irq
	wire         irq_mapper_receiver3_irq;                                   // uart_0:irq -> irq_mapper:receiver3_irq
	wire  [31:0] nios2_gen2_0_irq_irq;                                       // irq_mapper:sender_irq -> nios2_gen2_0:irq
	wire         rst_controller_reset_out_reset;                             // rst_controller:reset_out -> dma_rx_0:reset
	wire         nios2_gen2_0_debug_reset_request_reset;                     // nios2_gen2_0:debug_reset_request -> [rst_controller:reset_in1, rst_controller_001:reset_in1]
	wire         rst_controller_001_reset_out_reset;                         // rst_controller_001:reset_out -> [i_reg16_0:reset_n, i_reg16_1:reset_n, i_reg16_2:reset_n, i_reg16_3:reset_n, i_reg16_4:reset_n, i_reg16_5:reset_n, i_reg16_6:reset_n, i_reg32_0:reset_n, i_reg32_1:reset_n, i_reg32_2:reset_n, i_reg32_3:reset_n, i_reg32_4:reset_n, i_reg32_5:reset_n, i_reg32_6:reset_n, i_reg32_7:reset_n, mm_interconnect_0:dma_rx_0_reset_reset_bridge_in_reset_reset, mm_interconnect_0:timer_0_reset_reset_bridge_in_reset_reset, o_reg32_0:reset_n, o_reg32_10:reset_n, o_reg32_11:reset_n, o_reg32_12:reset_n, o_reg32_13:reset_n, o_reg32_1:reset_n, o_reg32_2:reset_n, o_reg32_3:reset_n, o_reg32_4:reset_n, o_reg32_5:reset_n, o_reg32_7:reset_n, o_reg32_8:reset_n, o_reg32_9:reset_n, timer_0:reset_n, timer_1:reset_n, uart_0:reset_n]
	wire         rst_controller_002_reset_out_reset;                         // rst_controller_002:reset_out -> [irq_mapper:reset, mm_interconnect_0:nios2_gen2_0_reset_reset_bridge_in_reset_reset, nios2_gen2_0:reset_n, o_reg32_6:reset_n, onchip_memory2_0:reset, rst_translator:in_reset]
	wire         rst_controller_002_reset_out_reset_req;                     // rst_controller_002:reset_req -> [nios2_gen2_0:reset_req, onchip_memory2_0:reset_req, rst_translator:reset_req_in]

	dma_receiver #(
		.DEPTH         (32),
		.clock_nsec    (20),
		.WATCHDOG_nsec (100000)
	) dma_rx_0 (
		.reset             (rst_controller_reset_out_reset),               //         reset.reset
		.av_mm_read        (mm_interconnect_0_dma_rx_0_av_mm_read),        //         av_mm.read
		.av_mm_readdata    (mm_interconnect_0_dma_rx_0_av_mm_readdata),    //              .readdata
		.av_mm_waitrequest (mm_interconnect_0_dma_rx_0_av_mm_waitrequest), //              .waitrequest
		.av_mm_write       (mm_interconnect_0_dma_rx_0_av_mm_write),       //              .write
		.av_mm_writedata   (mm_interconnect_0_dma_rx_0_av_mm_writedata),   //              .writedata
		.av_mm_addr        (mm_interconnect_0_dma_rx_0_av_mm_address),     //              .address
		.coe_RX_DONE       (coe_done),                                     // conduit_end_0.done
		.coe_RX_DATA       (coe_data),                                     //              .data
		.clock             (clk_clk)                                       //         clock.clk
	);

	NiosBase_i_reg16_0 i_reg16_0 (
		.clk      (clk_clk),                                 //                 clk.clk
		.reset_n  (~rst_controller_001_reset_out_reset),     //               reset.reset_n
		.address  (mm_interconnect_0_i_reg16_0_s1_address),  //                  s1.address
		.readdata (mm_interconnect_0_i_reg16_0_s1_readdata), //                    .readdata
		.in_port  (i_reg16_0_export)                         // external_connection.export
	);

	NiosBase_i_reg16_0 i_reg16_1 (
		.clk      (clk_clk),                                 //                 clk.clk
		.reset_n  (~rst_controller_001_reset_out_reset),     //               reset.reset_n
		.address  (mm_interconnect_0_i_reg16_1_s1_address),  //                  s1.address
		.readdata (mm_interconnect_0_i_reg16_1_s1_readdata), //                    .readdata
		.in_port  (i_reg16_1_export)                         // external_connection.export
	);

	NiosBase_i_reg16_0 i_reg16_2 (
		.clk      (clk_clk),                                 //                 clk.clk
		.reset_n  (~rst_controller_001_reset_out_reset),     //               reset.reset_n
		.address  (mm_interconnect_0_i_reg16_2_s1_address),  //                  s1.address
		.readdata (mm_interconnect_0_i_reg16_2_s1_readdata), //                    .readdata
		.in_port  (i_reg16_2_export)                         // external_connection.export
	);

	NiosBase_i_reg16_0 i_reg16_3 (
		.clk      (clk_clk),                                 //                 clk.clk
		.reset_n  (~rst_controller_001_reset_out_reset),     //               reset.reset_n
		.address  (mm_interconnect_0_i_reg16_3_s1_address),  //                  s1.address
		.readdata (mm_interconnect_0_i_reg16_3_s1_readdata), //                    .readdata
		.in_port  (i_reg16_3_export)                         // external_connection.export
	);

	NiosBase_i_reg16_0 i_reg16_4 (
		.clk      (clk_clk),                                 //                 clk.clk
		.reset_n  (~rst_controller_001_reset_out_reset),     //               reset.reset_n
		.address  (mm_interconnect_0_i_reg16_4_s1_address),  //                  s1.address
		.readdata (mm_interconnect_0_i_reg16_4_s1_readdata), //                    .readdata
		.in_port  (i_reg16_4_export)                         // external_connection.export
	);

	NiosBase_i_reg16_0 i_reg16_5 (
		.clk      (clk_clk),                                 //                 clk.clk
		.reset_n  (~rst_controller_001_reset_out_reset),     //               reset.reset_n
		.address  (mm_interconnect_0_i_reg16_5_s1_address),  //                  s1.address
		.readdata (mm_interconnect_0_i_reg16_5_s1_readdata), //                    .readdata
		.in_port  (i_reg16_5_export)                         // external_connection.export
	);

	NiosBase_i_reg16_0 i_reg16_6 (
		.clk      (clk_clk),                                 //                 clk.clk
		.reset_n  (~rst_controller_001_reset_out_reset),     //               reset.reset_n
		.address  (mm_interconnect_0_i_reg16_6_s1_address),  //                  s1.address
		.readdata (mm_interconnect_0_i_reg16_6_s1_readdata), //                    .readdata
		.in_port  (i_reg16_6_export)                         // external_connection.export
	);

	NiosBase_i_reg32_0 i_reg32_0 (
		.clk        (clk_clk),                                   //                 clk.clk
		.reset_n    (~rst_controller_001_reset_out_reset),       //               reset.reset_n
		.address    (mm_interconnect_0_i_reg32_0_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_i_reg32_0_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_i_reg32_0_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_i_reg32_0_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_i_reg32_0_s1_readdata),   //                    .readdata
		.in_port    (i_reg32_0_export),                          // external_connection.export
		.irq        (irq_mapper_receiver2_irq)                   //                 irq.irq
	);

	NiosBase_i_reg32_1 i_reg32_1 (
		.clk      (clk_clk),                                 //                 clk.clk
		.reset_n  (~rst_controller_001_reset_out_reset),     //               reset.reset_n
		.address  (mm_interconnect_0_i_reg32_1_s1_address),  //                  s1.address
		.readdata (mm_interconnect_0_i_reg32_1_s1_readdata), //                    .readdata
		.in_port  (i_reg32_1_export)                         // external_connection.export
	);

	NiosBase_i_reg32_1 i_reg32_2 (
		.clk      (clk_clk),                                 //                 clk.clk
		.reset_n  (~rst_controller_001_reset_out_reset),     //               reset.reset_n
		.address  (mm_interconnect_0_i_reg32_2_s1_address),  //                  s1.address
		.readdata (mm_interconnect_0_i_reg32_2_s1_readdata), //                    .readdata
		.in_port  (i_reg32_2_export)                         // external_connection.export
	);

	NiosBase_i_reg32_1 i_reg32_3 (
		.clk      (clk_clk),                                 //                 clk.clk
		.reset_n  (~rst_controller_001_reset_out_reset),     //               reset.reset_n
		.address  (mm_interconnect_0_i_reg32_3_s1_address),  //                  s1.address
		.readdata (mm_interconnect_0_i_reg32_3_s1_readdata), //                    .readdata
		.in_port  (i_reg32_3_export)                         // external_connection.export
	);

	NiosBase_i_reg32_1 i_reg32_4 (
		.clk      (clk_clk),                                 //                 clk.clk
		.reset_n  (~rst_controller_001_reset_out_reset),     //               reset.reset_n
		.address  (mm_interconnect_0_i_reg32_4_s1_address),  //                  s1.address
		.readdata (mm_interconnect_0_i_reg32_4_s1_readdata), //                    .readdata
		.in_port  (i_reg32_4_export)                         // external_connection.export
	);

	NiosBase_i_reg32_1 i_reg32_5 (
		.clk      (clk_clk),                                 //                 clk.clk
		.reset_n  (~rst_controller_001_reset_out_reset),     //               reset.reset_n
		.address  (mm_interconnect_0_i_reg32_5_s1_address),  //                  s1.address
		.readdata (mm_interconnect_0_i_reg32_5_s1_readdata), //                    .readdata
		.in_port  (i_reg32_5_export)                         // external_connection.export
	);

	NiosBase_i_reg32_1 i_reg32_6 (
		.clk      (clk_clk),                                 //                 clk.clk
		.reset_n  (~rst_controller_001_reset_out_reset),     //               reset.reset_n
		.address  (mm_interconnect_0_i_reg32_6_s1_address),  //                  s1.address
		.readdata (mm_interconnect_0_i_reg32_6_s1_readdata), //                    .readdata
		.in_port  (i_reg32_6_export)                         // external_connection.export
	);

	NiosBase_i_reg32_1 i_reg32_7 (
		.clk      (clk_clk),                                 //                 clk.clk
		.reset_n  (~rst_controller_001_reset_out_reset),     //               reset.reset_n
		.address  (mm_interconnect_0_i_reg32_7_s1_address),  //                  s1.address
		.readdata (mm_interconnect_0_i_reg32_7_s1_readdata), //                    .readdata
		.in_port  (i_reg32_7_export)                         // external_connection.export
	);

	NiosBase_nios2_gen2_0 nios2_gen2_0 (
		.clk                                 (clk_clk),                                                    //                       clk.clk
		.reset_n                             (~rst_controller_002_reset_out_reset),                        //                     reset.reset_n
		.reset_req                           (rst_controller_002_reset_out_reset_req),                     //                          .reset_req
		.d_address                           (nios2_gen2_0_data_master_address),                           //               data_master.address
		.d_byteenable                        (nios2_gen2_0_data_master_byteenable),                        //                          .byteenable
		.d_read                              (nios2_gen2_0_data_master_read),                              //                          .read
		.d_readdata                          (nios2_gen2_0_data_master_readdata),                          //                          .readdata
		.d_waitrequest                       (nios2_gen2_0_data_master_waitrequest),                       //                          .waitrequest
		.d_write                             (nios2_gen2_0_data_master_write),                             //                          .write
		.d_writedata                         (nios2_gen2_0_data_master_writedata),                         //                          .writedata
		.debug_mem_slave_debugaccess_to_roms (nios2_gen2_0_data_master_debugaccess),                       //                          .debugaccess
		.i_address                           (nios2_gen2_0_instruction_master_address),                    //        instruction_master.address
		.i_read                              (nios2_gen2_0_instruction_master_read),                       //                          .read
		.i_readdata                          (nios2_gen2_0_instruction_master_readdata),                   //                          .readdata
		.i_waitrequest                       (nios2_gen2_0_instruction_master_waitrequest),                //                          .waitrequest
		.irq                                 (nios2_gen2_0_irq_irq),                                       //                       irq.irq
		.debug_reset_request                 (nios2_gen2_0_debug_reset_request_reset),                     //       debug_reset_request.reset
		.debug_mem_slave_address             (mm_interconnect_0_nios2_gen2_0_debug_mem_slave_address),     //           debug_mem_slave.address
		.debug_mem_slave_byteenable          (mm_interconnect_0_nios2_gen2_0_debug_mem_slave_byteenable),  //                          .byteenable
		.debug_mem_slave_debugaccess         (mm_interconnect_0_nios2_gen2_0_debug_mem_slave_debugaccess), //                          .debugaccess
		.debug_mem_slave_read                (mm_interconnect_0_nios2_gen2_0_debug_mem_slave_read),        //                          .read
		.debug_mem_slave_readdata            (mm_interconnect_0_nios2_gen2_0_debug_mem_slave_readdata),    //                          .readdata
		.debug_mem_slave_waitrequest         (mm_interconnect_0_nios2_gen2_0_debug_mem_slave_waitrequest), //                          .waitrequest
		.debug_mem_slave_write               (mm_interconnect_0_nios2_gen2_0_debug_mem_slave_write),       //                          .write
		.debug_mem_slave_writedata           (mm_interconnect_0_nios2_gen2_0_debug_mem_slave_writedata),   //                          .writedata
		.dummy_ci_port                       ()                                                            // custom_instruction_master.readra
	);

	NiosBase_o_reg32_0 o_reg32_0 (
		.clk        (clk_clk),                                   //                 clk.clk
		.reset_n    (~rst_controller_001_reset_out_reset),       //               reset.reset_n
		.address    (mm_interconnect_0_o_reg32_0_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_o_reg32_0_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_o_reg32_0_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_o_reg32_0_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_o_reg32_0_s1_readdata),   //                    .readdata
		.out_port   (o_reg32_0_export)                           // external_connection.export
	);

	NiosBase_o_reg32_0 o_reg32_1 (
		.clk        (clk_clk),                                   //                 clk.clk
		.reset_n    (~rst_controller_001_reset_out_reset),       //               reset.reset_n
		.address    (mm_interconnect_0_o_reg32_1_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_o_reg32_1_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_o_reg32_1_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_o_reg32_1_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_o_reg32_1_s1_readdata),   //                    .readdata
		.out_port   (o_reg32_1_export)                           // external_connection.export
	);

	NiosBase_o_reg32_0 o_reg32_10 (
		.clk        (clk_clk),                                    //                 clk.clk
		.reset_n    (~rst_controller_001_reset_out_reset),        //               reset.reset_n
		.address    (mm_interconnect_0_o_reg32_10_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_o_reg32_10_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_o_reg32_10_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_o_reg32_10_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_o_reg32_10_s1_readdata),   //                    .readdata
		.out_port   (o_reg32_10_export)                           // external_connection.export
	);

	NiosBase_o_reg32_0 o_reg32_11 (
		.clk        (clk_clk),                                    //                 clk.clk
		.reset_n    (~rst_controller_001_reset_out_reset),        //               reset.reset_n
		.address    (mm_interconnect_0_o_reg32_11_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_o_reg32_11_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_o_reg32_11_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_o_reg32_11_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_o_reg32_11_s1_readdata),   //                    .readdata
		.out_port   (o_reg32_11_export)                           // external_connection.export
	);

	NiosBase_o_reg32_0 o_reg32_12 (
		.clk        (clk_clk),                                    //                 clk.clk
		.reset_n    (~rst_controller_001_reset_out_reset),        //               reset.reset_n
		.address    (mm_interconnect_0_o_reg32_12_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_o_reg32_12_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_o_reg32_12_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_o_reg32_12_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_o_reg32_12_s1_readdata),   //                    .readdata
		.out_port   (o_reg32_12_export)                           // external_connection.export
	);

	NiosBase_o_reg32_0 o_reg32_13 (
		.clk        (clk_clk),                                    //                 clk.clk
		.reset_n    (~rst_controller_001_reset_out_reset),        //               reset.reset_n
		.address    (mm_interconnect_0_o_reg32_13_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_o_reg32_13_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_o_reg32_13_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_o_reg32_13_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_o_reg32_13_s1_readdata),   //                    .readdata
		.out_port   (o_reg32_13_export)                           // external_connection.export
	);

	NiosBase_o_reg32_0 o_reg32_2 (
		.clk        (clk_clk),                                   //                 clk.clk
		.reset_n    (~rst_controller_001_reset_out_reset),       //               reset.reset_n
		.address    (mm_interconnect_0_o_reg32_2_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_o_reg32_2_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_o_reg32_2_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_o_reg32_2_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_o_reg32_2_s1_readdata),   //                    .readdata
		.out_port   (o_reg32_2_export)                           // external_connection.export
	);

	NiosBase_o_reg32_0 o_reg32_3 (
		.clk        (clk_clk),                                   //                 clk.clk
		.reset_n    (~rst_controller_001_reset_out_reset),       //               reset.reset_n
		.address    (mm_interconnect_0_o_reg32_3_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_o_reg32_3_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_o_reg32_3_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_o_reg32_3_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_o_reg32_3_s1_readdata),   //                    .readdata
		.out_port   (o_reg32_3_export)                           // external_connection.export
	);

	NiosBase_o_reg32_0 o_reg32_4 (
		.clk        (clk_clk),                                   //                 clk.clk
		.reset_n    (~rst_controller_001_reset_out_reset),       //               reset.reset_n
		.address    (mm_interconnect_0_o_reg32_4_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_o_reg32_4_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_o_reg32_4_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_o_reg32_4_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_o_reg32_4_s1_readdata),   //                    .readdata
		.out_port   (o_reg32_4_export)                           // external_connection.export
	);

	NiosBase_o_reg32_0 o_reg32_5 (
		.clk        (clk_clk),                                   //                 clk.clk
		.reset_n    (~rst_controller_001_reset_out_reset),       //               reset.reset_n
		.address    (mm_interconnect_0_o_reg32_5_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_o_reg32_5_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_o_reg32_5_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_o_reg32_5_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_o_reg32_5_s1_readdata),   //                    .readdata
		.out_port   (o_reg32_5_export)                           // external_connection.export
	);

	NiosBase_o_reg32_0 o_reg32_6 (
		.clk        (clk_clk),                                   //                 clk.clk
		.reset_n    (~rst_controller_002_reset_out_reset),       //               reset.reset_n
		.address    (mm_interconnect_0_o_reg32_6_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_o_reg32_6_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_o_reg32_6_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_o_reg32_6_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_o_reg32_6_s1_readdata),   //                    .readdata
		.out_port   (o_reg32_6_export)                           // external_connection.export
	);

	NiosBase_o_reg32_0 o_reg32_7 (
		.clk        (clk_clk),                                   //                 clk.clk
		.reset_n    (~rst_controller_001_reset_out_reset),       //               reset.reset_n
		.address    (mm_interconnect_0_o_reg32_7_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_o_reg32_7_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_o_reg32_7_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_o_reg32_7_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_o_reg32_7_s1_readdata),   //                    .readdata
		.out_port   (o_reg32_7_export)                           // external_connection.export
	);

	NiosBase_o_reg32_0 o_reg32_8 (
		.clk        (clk_clk),                                   //                 clk.clk
		.reset_n    (~rst_controller_001_reset_out_reset),       //               reset.reset_n
		.address    (mm_interconnect_0_o_reg32_8_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_o_reg32_8_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_o_reg32_8_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_o_reg32_8_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_o_reg32_8_s1_readdata),   //                    .readdata
		.out_port   (o_reg32_8_export)                           // external_connection.export
	);

	NiosBase_o_reg32_0 o_reg32_9 (
		.clk        (clk_clk),                                   //                 clk.clk
		.reset_n    (~rst_controller_001_reset_out_reset),       //               reset.reset_n
		.address    (mm_interconnect_0_o_reg32_9_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_o_reg32_9_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_o_reg32_9_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_o_reg32_9_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_o_reg32_9_s1_readdata),   //                    .readdata
		.out_port   (o_reg32_9_export)                           // external_connection.export
	);

	NiosBase_onchip_memory2_0 onchip_memory2_0 (
		.clk        (clk_clk),                                          //   clk1.clk
		.address    (mm_interconnect_0_onchip_memory2_0_s1_address),    //     s1.address
		.clken      (mm_interconnect_0_onchip_memory2_0_s1_clken),      //       .clken
		.chipselect (mm_interconnect_0_onchip_memory2_0_s1_chipselect), //       .chipselect
		.write      (mm_interconnect_0_onchip_memory2_0_s1_write),      //       .write
		.readdata   (mm_interconnect_0_onchip_memory2_0_s1_readdata),   //       .readdata
		.writedata  (mm_interconnect_0_onchip_memory2_0_s1_writedata),  //       .writedata
		.byteenable (mm_interconnect_0_onchip_memory2_0_s1_byteenable), //       .byteenable
		.reset      (rst_controller_002_reset_out_reset),               // reset1.reset
		.reset_req  (rst_controller_002_reset_out_reset_req),           //       .reset_req
		.freeze     (1'b0)                                              // (terminated)
	);

	NiosBase_timer_0 timer_0 (
		.clk        (clk_clk),                                 //   clk.clk
		.reset_n    (~rst_controller_001_reset_out_reset),     // reset.reset_n
		.address    (mm_interconnect_0_timer_0_s1_address),    //    s1.address
		.writedata  (mm_interconnect_0_timer_0_s1_writedata),  //      .writedata
		.readdata   (mm_interconnect_0_timer_0_s1_readdata),   //      .readdata
		.chipselect (mm_interconnect_0_timer_0_s1_chipselect), //      .chipselect
		.write_n    (~mm_interconnect_0_timer_0_s1_write),     //      .write_n
		.irq        (irq_mapper_receiver0_irq)                 //   irq.irq
	);

	NiosBase_timer_1 timer_1 (
		.clk        (clk_clk),                                 //   clk.clk
		.reset_n    (~rst_controller_001_reset_out_reset),     // reset.reset_n
		.address    (mm_interconnect_0_timer_1_s1_address),    //    s1.address
		.writedata  (mm_interconnect_0_timer_1_s1_writedata),  //      .writedata
		.readdata   (mm_interconnect_0_timer_1_s1_readdata),   //      .readdata
		.chipselect (mm_interconnect_0_timer_1_s1_chipselect), //      .chipselect
		.write_n    (~mm_interconnect_0_timer_1_s1_write),     //      .write_n
		.irq        (irq_mapper_receiver1_irq)                 //   irq.irq
	);

	NiosBase_uart_0 uart_0 (
		.clk           (clk_clk),                                   //                 clk.clk
		.reset_n       (~rst_controller_001_reset_out_reset),       //               reset.reset_n
		.address       (mm_interconnect_0_uart_0_s1_address),       //                  s1.address
		.begintransfer (mm_interconnect_0_uart_0_s1_begintransfer), //                    .begintransfer
		.chipselect    (mm_interconnect_0_uart_0_s1_chipselect),    //                    .chipselect
		.read_n        (~mm_interconnect_0_uart_0_s1_read),         //                    .read_n
		.write_n       (~mm_interconnect_0_uart_0_s1_write),        //                    .write_n
		.writedata     (mm_interconnect_0_uart_0_s1_writedata),     //                    .writedata
		.readdata      (mm_interconnect_0_uart_0_s1_readdata),      //                    .readdata
		.rxd           (uart_rxd),                                  // external_connection.export
		.txd           (uart_txd),                                  //                    .export
		.irq           (irq_mapper_receiver3_irq)                   //                 irq.irq
	);

	NiosBase_mm_interconnect_0 mm_interconnect_0 (
		.clk_0_clk_clk                                  (clk_clk),                                                    //                                clk_0_clk.clk
		.dma_rx_0_reset_reset_bridge_in_reset_reset     (rst_controller_001_reset_out_reset),                         //     dma_rx_0_reset_reset_bridge_in_reset.reset
		.nios2_gen2_0_reset_reset_bridge_in_reset_reset (rst_controller_002_reset_out_reset),                         // nios2_gen2_0_reset_reset_bridge_in_reset.reset
		.timer_0_reset_reset_bridge_in_reset_reset      (rst_controller_001_reset_out_reset),                         //      timer_0_reset_reset_bridge_in_reset.reset
		.nios2_gen2_0_data_master_address               (nios2_gen2_0_data_master_address),                           //                 nios2_gen2_0_data_master.address
		.nios2_gen2_0_data_master_waitrequest           (nios2_gen2_0_data_master_waitrequest),                       //                                         .waitrequest
		.nios2_gen2_0_data_master_byteenable            (nios2_gen2_0_data_master_byteenable),                        //                                         .byteenable
		.nios2_gen2_0_data_master_read                  (nios2_gen2_0_data_master_read),                              //                                         .read
		.nios2_gen2_0_data_master_readdata              (nios2_gen2_0_data_master_readdata),                          //                                         .readdata
		.nios2_gen2_0_data_master_write                 (nios2_gen2_0_data_master_write),                             //                                         .write
		.nios2_gen2_0_data_master_writedata             (nios2_gen2_0_data_master_writedata),                         //                                         .writedata
		.nios2_gen2_0_data_master_debugaccess           (nios2_gen2_0_data_master_debugaccess),                       //                                         .debugaccess
		.nios2_gen2_0_instruction_master_address        (nios2_gen2_0_instruction_master_address),                    //          nios2_gen2_0_instruction_master.address
		.nios2_gen2_0_instruction_master_waitrequest    (nios2_gen2_0_instruction_master_waitrequest),                //                                         .waitrequest
		.nios2_gen2_0_instruction_master_read           (nios2_gen2_0_instruction_master_read),                       //                                         .read
		.nios2_gen2_0_instruction_master_readdata       (nios2_gen2_0_instruction_master_readdata),                   //                                         .readdata
		.dma_rx_0_av_mm_address                         (mm_interconnect_0_dma_rx_0_av_mm_address),                   //                           dma_rx_0_av_mm.address
		.dma_rx_0_av_mm_write                           (mm_interconnect_0_dma_rx_0_av_mm_write),                     //                                         .write
		.dma_rx_0_av_mm_read                            (mm_interconnect_0_dma_rx_0_av_mm_read),                      //                                         .read
		.dma_rx_0_av_mm_readdata                        (mm_interconnect_0_dma_rx_0_av_mm_readdata),                  //                                         .readdata
		.dma_rx_0_av_mm_writedata                       (mm_interconnect_0_dma_rx_0_av_mm_writedata),                 //                                         .writedata
		.dma_rx_0_av_mm_waitrequest                     (mm_interconnect_0_dma_rx_0_av_mm_waitrequest),               //                                         .waitrequest
		.i_reg16_0_s1_address                           (mm_interconnect_0_i_reg16_0_s1_address),                     //                             i_reg16_0_s1.address
		.i_reg16_0_s1_readdata                          (mm_interconnect_0_i_reg16_0_s1_readdata),                    //                                         .readdata
		.i_reg16_1_s1_address                           (mm_interconnect_0_i_reg16_1_s1_address),                     //                             i_reg16_1_s1.address
		.i_reg16_1_s1_readdata                          (mm_interconnect_0_i_reg16_1_s1_readdata),                    //                                         .readdata
		.i_reg16_2_s1_address                           (mm_interconnect_0_i_reg16_2_s1_address),                     //                             i_reg16_2_s1.address
		.i_reg16_2_s1_readdata                          (mm_interconnect_0_i_reg16_2_s1_readdata),                    //                                         .readdata
		.i_reg16_3_s1_address                           (mm_interconnect_0_i_reg16_3_s1_address),                     //                             i_reg16_3_s1.address
		.i_reg16_3_s1_readdata                          (mm_interconnect_0_i_reg16_3_s1_readdata),                    //                                         .readdata
		.i_reg16_4_s1_address                           (mm_interconnect_0_i_reg16_4_s1_address),                     //                             i_reg16_4_s1.address
		.i_reg16_4_s1_readdata                          (mm_interconnect_0_i_reg16_4_s1_readdata),                    //                                         .readdata
		.i_reg16_5_s1_address                           (mm_interconnect_0_i_reg16_5_s1_address),                     //                             i_reg16_5_s1.address
		.i_reg16_5_s1_readdata                          (mm_interconnect_0_i_reg16_5_s1_readdata),                    //                                         .readdata
		.i_reg16_6_s1_address                           (mm_interconnect_0_i_reg16_6_s1_address),                     //                             i_reg16_6_s1.address
		.i_reg16_6_s1_readdata                          (mm_interconnect_0_i_reg16_6_s1_readdata),                    //                                         .readdata
		.i_reg32_0_s1_address                           (mm_interconnect_0_i_reg32_0_s1_address),                     //                             i_reg32_0_s1.address
		.i_reg32_0_s1_write                             (mm_interconnect_0_i_reg32_0_s1_write),                       //                                         .write
		.i_reg32_0_s1_readdata                          (mm_interconnect_0_i_reg32_0_s1_readdata),                    //                                         .readdata
		.i_reg32_0_s1_writedata                         (mm_interconnect_0_i_reg32_0_s1_writedata),                   //                                         .writedata
		.i_reg32_0_s1_chipselect                        (mm_interconnect_0_i_reg32_0_s1_chipselect),                  //                                         .chipselect
		.i_reg32_1_s1_address                           (mm_interconnect_0_i_reg32_1_s1_address),                     //                             i_reg32_1_s1.address
		.i_reg32_1_s1_readdata                          (mm_interconnect_0_i_reg32_1_s1_readdata),                    //                                         .readdata
		.i_reg32_2_s1_address                           (mm_interconnect_0_i_reg32_2_s1_address),                     //                             i_reg32_2_s1.address
		.i_reg32_2_s1_readdata                          (mm_interconnect_0_i_reg32_2_s1_readdata),                    //                                         .readdata
		.i_reg32_3_s1_address                           (mm_interconnect_0_i_reg32_3_s1_address),                     //                             i_reg32_3_s1.address
		.i_reg32_3_s1_readdata                          (mm_interconnect_0_i_reg32_3_s1_readdata),                    //                                         .readdata
		.i_reg32_4_s1_address                           (mm_interconnect_0_i_reg32_4_s1_address),                     //                             i_reg32_4_s1.address
		.i_reg32_4_s1_readdata                          (mm_interconnect_0_i_reg32_4_s1_readdata),                    //                                         .readdata
		.i_reg32_5_s1_address                           (mm_interconnect_0_i_reg32_5_s1_address),                     //                             i_reg32_5_s1.address
		.i_reg32_5_s1_readdata                          (mm_interconnect_0_i_reg32_5_s1_readdata),                    //                                         .readdata
		.i_reg32_6_s1_address                           (mm_interconnect_0_i_reg32_6_s1_address),                     //                             i_reg32_6_s1.address
		.i_reg32_6_s1_readdata                          (mm_interconnect_0_i_reg32_6_s1_readdata),                    //                                         .readdata
		.i_reg32_7_s1_address                           (mm_interconnect_0_i_reg32_7_s1_address),                     //                             i_reg32_7_s1.address
		.i_reg32_7_s1_readdata                          (mm_interconnect_0_i_reg32_7_s1_readdata),                    //                                         .readdata
		.nios2_gen2_0_debug_mem_slave_address           (mm_interconnect_0_nios2_gen2_0_debug_mem_slave_address),     //             nios2_gen2_0_debug_mem_slave.address
		.nios2_gen2_0_debug_mem_slave_write             (mm_interconnect_0_nios2_gen2_0_debug_mem_slave_write),       //                                         .write
		.nios2_gen2_0_debug_mem_slave_read              (mm_interconnect_0_nios2_gen2_0_debug_mem_slave_read),        //                                         .read
		.nios2_gen2_0_debug_mem_slave_readdata          (mm_interconnect_0_nios2_gen2_0_debug_mem_slave_readdata),    //                                         .readdata
		.nios2_gen2_0_debug_mem_slave_writedata         (mm_interconnect_0_nios2_gen2_0_debug_mem_slave_writedata),   //                                         .writedata
		.nios2_gen2_0_debug_mem_slave_byteenable        (mm_interconnect_0_nios2_gen2_0_debug_mem_slave_byteenable),  //                                         .byteenable
		.nios2_gen2_0_debug_mem_slave_waitrequest       (mm_interconnect_0_nios2_gen2_0_debug_mem_slave_waitrequest), //                                         .waitrequest
		.nios2_gen2_0_debug_mem_slave_debugaccess       (mm_interconnect_0_nios2_gen2_0_debug_mem_slave_debugaccess), //                                         .debugaccess
		.o_reg32_0_s1_address                           (mm_interconnect_0_o_reg32_0_s1_address),                     //                             o_reg32_0_s1.address
		.o_reg32_0_s1_write                             (mm_interconnect_0_o_reg32_0_s1_write),                       //                                         .write
		.o_reg32_0_s1_readdata                          (mm_interconnect_0_o_reg32_0_s1_readdata),                    //                                         .readdata
		.o_reg32_0_s1_writedata                         (mm_interconnect_0_o_reg32_0_s1_writedata),                   //                                         .writedata
		.o_reg32_0_s1_chipselect                        (mm_interconnect_0_o_reg32_0_s1_chipselect),                  //                                         .chipselect
		.o_reg32_1_s1_address                           (mm_interconnect_0_o_reg32_1_s1_address),                     //                             o_reg32_1_s1.address
		.o_reg32_1_s1_write                             (mm_interconnect_0_o_reg32_1_s1_write),                       //                                         .write
		.o_reg32_1_s1_readdata                          (mm_interconnect_0_o_reg32_1_s1_readdata),                    //                                         .readdata
		.o_reg32_1_s1_writedata                         (mm_interconnect_0_o_reg32_1_s1_writedata),                   //                                         .writedata
		.o_reg32_1_s1_chipselect                        (mm_interconnect_0_o_reg32_1_s1_chipselect),                  //                                         .chipselect
		.o_reg32_10_s1_address                          (mm_interconnect_0_o_reg32_10_s1_address),                    //                            o_reg32_10_s1.address
		.o_reg32_10_s1_write                            (mm_interconnect_0_o_reg32_10_s1_write),                      //                                         .write
		.o_reg32_10_s1_readdata                         (mm_interconnect_0_o_reg32_10_s1_readdata),                   //                                         .readdata
		.o_reg32_10_s1_writedata                        (mm_interconnect_0_o_reg32_10_s1_writedata),                  //                                         .writedata
		.o_reg32_10_s1_chipselect                       (mm_interconnect_0_o_reg32_10_s1_chipselect),                 //                                         .chipselect
		.o_reg32_11_s1_address                          (mm_interconnect_0_o_reg32_11_s1_address),                    //                            o_reg32_11_s1.address
		.o_reg32_11_s1_write                            (mm_interconnect_0_o_reg32_11_s1_write),                      //                                         .write
		.o_reg32_11_s1_readdata                         (mm_interconnect_0_o_reg32_11_s1_readdata),                   //                                         .readdata
		.o_reg32_11_s1_writedata                        (mm_interconnect_0_o_reg32_11_s1_writedata),                  //                                         .writedata
		.o_reg32_11_s1_chipselect                       (mm_interconnect_0_o_reg32_11_s1_chipselect),                 //                                         .chipselect
		.o_reg32_12_s1_address                          (mm_interconnect_0_o_reg32_12_s1_address),                    //                            o_reg32_12_s1.address
		.o_reg32_12_s1_write                            (mm_interconnect_0_o_reg32_12_s1_write),                      //                                         .write
		.o_reg32_12_s1_readdata                         (mm_interconnect_0_o_reg32_12_s1_readdata),                   //                                         .readdata
		.o_reg32_12_s1_writedata                        (mm_interconnect_0_o_reg32_12_s1_writedata),                  //                                         .writedata
		.o_reg32_12_s1_chipselect                       (mm_interconnect_0_o_reg32_12_s1_chipselect),                 //                                         .chipselect
		.o_reg32_13_s1_address                          (mm_interconnect_0_o_reg32_13_s1_address),                    //                            o_reg32_13_s1.address
		.o_reg32_13_s1_write                            (mm_interconnect_0_o_reg32_13_s1_write),                      //                                         .write
		.o_reg32_13_s1_readdata                         (mm_interconnect_0_o_reg32_13_s1_readdata),                   //                                         .readdata
		.o_reg32_13_s1_writedata                        (mm_interconnect_0_o_reg32_13_s1_writedata),                  //                                         .writedata
		.o_reg32_13_s1_chipselect                       (mm_interconnect_0_o_reg32_13_s1_chipselect),                 //                                         .chipselect
		.o_reg32_2_s1_address                           (mm_interconnect_0_o_reg32_2_s1_address),                     //                             o_reg32_2_s1.address
		.o_reg32_2_s1_write                             (mm_interconnect_0_o_reg32_2_s1_write),                       //                                         .write
		.o_reg32_2_s1_readdata                          (mm_interconnect_0_o_reg32_2_s1_readdata),                    //                                         .readdata
		.o_reg32_2_s1_writedata                         (mm_interconnect_0_o_reg32_2_s1_writedata),                   //                                         .writedata
		.o_reg32_2_s1_chipselect                        (mm_interconnect_0_o_reg32_2_s1_chipselect),                  //                                         .chipselect
		.o_reg32_3_s1_address                           (mm_interconnect_0_o_reg32_3_s1_address),                     //                             o_reg32_3_s1.address
		.o_reg32_3_s1_write                             (mm_interconnect_0_o_reg32_3_s1_write),                       //                                         .write
		.o_reg32_3_s1_readdata                          (mm_interconnect_0_o_reg32_3_s1_readdata),                    //                                         .readdata
		.o_reg32_3_s1_writedata                         (mm_interconnect_0_o_reg32_3_s1_writedata),                   //                                         .writedata
		.o_reg32_3_s1_chipselect                        (mm_interconnect_0_o_reg32_3_s1_chipselect),                  //                                         .chipselect
		.o_reg32_4_s1_address                           (mm_interconnect_0_o_reg32_4_s1_address),                     //                             o_reg32_4_s1.address
		.o_reg32_4_s1_write                             (mm_interconnect_0_o_reg32_4_s1_write),                       //                                         .write
		.o_reg32_4_s1_readdata                          (mm_interconnect_0_o_reg32_4_s1_readdata),                    //                                         .readdata
		.o_reg32_4_s1_writedata                         (mm_interconnect_0_o_reg32_4_s1_writedata),                   //                                         .writedata
		.o_reg32_4_s1_chipselect                        (mm_interconnect_0_o_reg32_4_s1_chipselect),                  //                                         .chipselect
		.o_reg32_5_s1_address                           (mm_interconnect_0_o_reg32_5_s1_address),                     //                             o_reg32_5_s1.address
		.o_reg32_5_s1_write                             (mm_interconnect_0_o_reg32_5_s1_write),                       //                                         .write
		.o_reg32_5_s1_readdata                          (mm_interconnect_0_o_reg32_5_s1_readdata),                    //                                         .readdata
		.o_reg32_5_s1_writedata                         (mm_interconnect_0_o_reg32_5_s1_writedata),                   //                                         .writedata
		.o_reg32_5_s1_chipselect                        (mm_interconnect_0_o_reg32_5_s1_chipselect),                  //                                         .chipselect
		.o_reg32_6_s1_address                           (mm_interconnect_0_o_reg32_6_s1_address),                     //                             o_reg32_6_s1.address
		.o_reg32_6_s1_write                             (mm_interconnect_0_o_reg32_6_s1_write),                       //                                         .write
		.o_reg32_6_s1_readdata                          (mm_interconnect_0_o_reg32_6_s1_readdata),                    //                                         .readdata
		.o_reg32_6_s1_writedata                         (mm_interconnect_0_o_reg32_6_s1_writedata),                   //                                         .writedata
		.o_reg32_6_s1_chipselect                        (mm_interconnect_0_o_reg32_6_s1_chipselect),                  //                                         .chipselect
		.o_reg32_7_s1_address                           (mm_interconnect_0_o_reg32_7_s1_address),                     //                             o_reg32_7_s1.address
		.o_reg32_7_s1_write                             (mm_interconnect_0_o_reg32_7_s1_write),                       //                                         .write
		.o_reg32_7_s1_readdata                          (mm_interconnect_0_o_reg32_7_s1_readdata),                    //                                         .readdata
		.o_reg32_7_s1_writedata                         (mm_interconnect_0_o_reg32_7_s1_writedata),                   //                                         .writedata
		.o_reg32_7_s1_chipselect                        (mm_interconnect_0_o_reg32_7_s1_chipselect),                  //                                         .chipselect
		.o_reg32_8_s1_address                           (mm_interconnect_0_o_reg32_8_s1_address),                     //                             o_reg32_8_s1.address
		.o_reg32_8_s1_write                             (mm_interconnect_0_o_reg32_8_s1_write),                       //                                         .write
		.o_reg32_8_s1_readdata                          (mm_interconnect_0_o_reg32_8_s1_readdata),                    //                                         .readdata
		.o_reg32_8_s1_writedata                         (mm_interconnect_0_o_reg32_8_s1_writedata),                   //                                         .writedata
		.o_reg32_8_s1_chipselect                        (mm_interconnect_0_o_reg32_8_s1_chipselect),                  //                                         .chipselect
		.o_reg32_9_s1_address                           (mm_interconnect_0_o_reg32_9_s1_address),                     //                             o_reg32_9_s1.address
		.o_reg32_9_s1_write                             (mm_interconnect_0_o_reg32_9_s1_write),                       //                                         .write
		.o_reg32_9_s1_readdata                          (mm_interconnect_0_o_reg32_9_s1_readdata),                    //                                         .readdata
		.o_reg32_9_s1_writedata                         (mm_interconnect_0_o_reg32_9_s1_writedata),                   //                                         .writedata
		.o_reg32_9_s1_chipselect                        (mm_interconnect_0_o_reg32_9_s1_chipselect),                  //                                         .chipselect
		.onchip_memory2_0_s1_address                    (mm_interconnect_0_onchip_memory2_0_s1_address),              //                      onchip_memory2_0_s1.address
		.onchip_memory2_0_s1_write                      (mm_interconnect_0_onchip_memory2_0_s1_write),                //                                         .write
		.onchip_memory2_0_s1_readdata                   (mm_interconnect_0_onchip_memory2_0_s1_readdata),             //                                         .readdata
		.onchip_memory2_0_s1_writedata                  (mm_interconnect_0_onchip_memory2_0_s1_writedata),            //                                         .writedata
		.onchip_memory2_0_s1_byteenable                 (mm_interconnect_0_onchip_memory2_0_s1_byteenable),           //                                         .byteenable
		.onchip_memory2_0_s1_chipselect                 (mm_interconnect_0_onchip_memory2_0_s1_chipselect),           //                                         .chipselect
		.onchip_memory2_0_s1_clken                      (mm_interconnect_0_onchip_memory2_0_s1_clken),                //                                         .clken
		.timer_0_s1_address                             (mm_interconnect_0_timer_0_s1_address),                       //                               timer_0_s1.address
		.timer_0_s1_write                               (mm_interconnect_0_timer_0_s1_write),                         //                                         .write
		.timer_0_s1_readdata                            (mm_interconnect_0_timer_0_s1_readdata),                      //                                         .readdata
		.timer_0_s1_writedata                           (mm_interconnect_0_timer_0_s1_writedata),                     //                                         .writedata
		.timer_0_s1_chipselect                          (mm_interconnect_0_timer_0_s1_chipselect),                    //                                         .chipselect
		.timer_1_s1_address                             (mm_interconnect_0_timer_1_s1_address),                       //                               timer_1_s1.address
		.timer_1_s1_write                               (mm_interconnect_0_timer_1_s1_write),                         //                                         .write
		.timer_1_s1_readdata                            (mm_interconnect_0_timer_1_s1_readdata),                      //                                         .readdata
		.timer_1_s1_writedata                           (mm_interconnect_0_timer_1_s1_writedata),                     //                                         .writedata
		.timer_1_s1_chipselect                          (mm_interconnect_0_timer_1_s1_chipselect),                    //                                         .chipselect
		.uart_0_s1_address                              (mm_interconnect_0_uart_0_s1_address),                        //                                uart_0_s1.address
		.uart_0_s1_write                                (mm_interconnect_0_uart_0_s1_write),                          //                                         .write
		.uart_0_s1_read                                 (mm_interconnect_0_uart_0_s1_read),                           //                                         .read
		.uart_0_s1_readdata                             (mm_interconnect_0_uart_0_s1_readdata),                       //                                         .readdata
		.uart_0_s1_writedata                            (mm_interconnect_0_uart_0_s1_writedata),                      //                                         .writedata
		.uart_0_s1_begintransfer                        (mm_interconnect_0_uart_0_s1_begintransfer),                  //                                         .begintransfer
		.uart_0_s1_chipselect                           (mm_interconnect_0_uart_0_s1_chipselect)                      //                                         .chipselect
	);

	NiosBase_irq_mapper irq_mapper (
		.clk           (clk_clk),                            //       clk.clk
		.reset         (rst_controller_002_reset_out_reset), // clk_reset.reset
		.receiver0_irq (irq_mapper_receiver0_irq),           // receiver0.irq
		.receiver1_irq (irq_mapper_receiver1_irq),           // receiver1.irq
		.receiver2_irq (irq_mapper_receiver2_irq),           // receiver2.irq
		.receiver3_irq (irq_mapper_receiver3_irq),           // receiver3.irq
		.sender_irq    (nios2_gen2_0_irq_irq)                //    sender.irq
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS          (2),
		.OUTPUT_RESET_SYNC_EDGES   ("both"),
		.SYNC_DEPTH                (2),
		.RESET_REQUEST_PRESENT     (0),
		.RESET_REQ_WAIT_TIME       (1),
		.MIN_RST_ASSERTION_TIME    (3),
		.RESET_REQ_EARLY_DSRT_TIME (1),
		.USE_RESET_REQUEST_IN0     (0),
		.USE_RESET_REQUEST_IN1     (0),
		.USE_RESET_REQUEST_IN2     (0),
		.USE_RESET_REQUEST_IN3     (0),
		.USE_RESET_REQUEST_IN4     (0),
		.USE_RESET_REQUEST_IN5     (0),
		.USE_RESET_REQUEST_IN6     (0),
		.USE_RESET_REQUEST_IN7     (0),
		.USE_RESET_REQUEST_IN8     (0),
		.USE_RESET_REQUEST_IN9     (0),
		.USE_RESET_REQUEST_IN10    (0),
		.USE_RESET_REQUEST_IN11    (0),
		.USE_RESET_REQUEST_IN12    (0),
		.USE_RESET_REQUEST_IN13    (0),
		.USE_RESET_REQUEST_IN14    (0),
		.USE_RESET_REQUEST_IN15    (0),
		.ADAPT_RESET_REQUEST       (0)
	) rst_controller (
		.reset_in0      (~reset_reset_n),                         // reset_in0.reset
		.reset_in1      (nios2_gen2_0_debug_reset_request_reset), // reset_in1.reset
		.clk            (clk_clk),                                //       clk.clk
		.reset_out      (rst_controller_reset_out_reset),         // reset_out.reset
		.reset_req      (),                                       // (terminated)
		.reset_req_in0  (1'b0),                                   // (terminated)
		.reset_req_in1  (1'b0),                                   // (terminated)
		.reset_in2      (1'b0),                                   // (terminated)
		.reset_req_in2  (1'b0),                                   // (terminated)
		.reset_in3      (1'b0),                                   // (terminated)
		.reset_req_in3  (1'b0),                                   // (terminated)
		.reset_in4      (1'b0),                                   // (terminated)
		.reset_req_in4  (1'b0),                                   // (terminated)
		.reset_in5      (1'b0),                                   // (terminated)
		.reset_req_in5  (1'b0),                                   // (terminated)
		.reset_in6      (1'b0),                                   // (terminated)
		.reset_req_in6  (1'b0),                                   // (terminated)
		.reset_in7      (1'b0),                                   // (terminated)
		.reset_req_in7  (1'b0),                                   // (terminated)
		.reset_in8      (1'b0),                                   // (terminated)
		.reset_req_in8  (1'b0),                                   // (terminated)
		.reset_in9      (1'b0),                                   // (terminated)
		.reset_req_in9  (1'b0),                                   // (terminated)
		.reset_in10     (1'b0),                                   // (terminated)
		.reset_req_in10 (1'b0),                                   // (terminated)
		.reset_in11     (1'b0),                                   // (terminated)
		.reset_req_in11 (1'b0),                                   // (terminated)
		.reset_in12     (1'b0),                                   // (terminated)
		.reset_req_in12 (1'b0),                                   // (terminated)
		.reset_in13     (1'b0),                                   // (terminated)
		.reset_req_in13 (1'b0),                                   // (terminated)
		.reset_in14     (1'b0),                                   // (terminated)
		.reset_req_in14 (1'b0),                                   // (terminated)
		.reset_in15     (1'b0),                                   // (terminated)
		.reset_req_in15 (1'b0)                                    // (terminated)
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS          (2),
		.OUTPUT_RESET_SYNC_EDGES   ("deassert"),
		.SYNC_DEPTH                (2),
		.RESET_REQUEST_PRESENT     (0),
		.RESET_REQ_WAIT_TIME       (1),
		.MIN_RST_ASSERTION_TIME    (3),
		.RESET_REQ_EARLY_DSRT_TIME (1),
		.USE_RESET_REQUEST_IN0     (0),
		.USE_RESET_REQUEST_IN1     (0),
		.USE_RESET_REQUEST_IN2     (0),
		.USE_RESET_REQUEST_IN3     (0),
		.USE_RESET_REQUEST_IN4     (0),
		.USE_RESET_REQUEST_IN5     (0),
		.USE_RESET_REQUEST_IN6     (0),
		.USE_RESET_REQUEST_IN7     (0),
		.USE_RESET_REQUEST_IN8     (0),
		.USE_RESET_REQUEST_IN9     (0),
		.USE_RESET_REQUEST_IN10    (0),
		.USE_RESET_REQUEST_IN11    (0),
		.USE_RESET_REQUEST_IN12    (0),
		.USE_RESET_REQUEST_IN13    (0),
		.USE_RESET_REQUEST_IN14    (0),
		.USE_RESET_REQUEST_IN15    (0),
		.ADAPT_RESET_REQUEST       (0)
	) rst_controller_001 (
		.reset_in0      (~reset_reset_n),                         // reset_in0.reset
		.reset_in1      (nios2_gen2_0_debug_reset_request_reset), // reset_in1.reset
		.clk            (clk_clk),                                //       clk.clk
		.reset_out      (rst_controller_001_reset_out_reset),     // reset_out.reset
		.reset_req      (),                                       // (terminated)
		.reset_req_in0  (1'b0),                                   // (terminated)
		.reset_req_in1  (1'b0),                                   // (terminated)
		.reset_in2      (1'b0),                                   // (terminated)
		.reset_req_in2  (1'b0),                                   // (terminated)
		.reset_in3      (1'b0),                                   // (terminated)
		.reset_req_in3  (1'b0),                                   // (terminated)
		.reset_in4      (1'b0),                                   // (terminated)
		.reset_req_in4  (1'b0),                                   // (terminated)
		.reset_in5      (1'b0),                                   // (terminated)
		.reset_req_in5  (1'b0),                                   // (terminated)
		.reset_in6      (1'b0),                                   // (terminated)
		.reset_req_in6  (1'b0),                                   // (terminated)
		.reset_in7      (1'b0),                                   // (terminated)
		.reset_req_in7  (1'b0),                                   // (terminated)
		.reset_in8      (1'b0),                                   // (terminated)
		.reset_req_in8  (1'b0),                                   // (terminated)
		.reset_in9      (1'b0),                                   // (terminated)
		.reset_req_in9  (1'b0),                                   // (terminated)
		.reset_in10     (1'b0),                                   // (terminated)
		.reset_req_in10 (1'b0),                                   // (terminated)
		.reset_in11     (1'b0),                                   // (terminated)
		.reset_req_in11 (1'b0),                                   // (terminated)
		.reset_in12     (1'b0),                                   // (terminated)
		.reset_req_in12 (1'b0),                                   // (terminated)
		.reset_in13     (1'b0),                                   // (terminated)
		.reset_req_in13 (1'b0),                                   // (terminated)
		.reset_in14     (1'b0),                                   // (terminated)
		.reset_req_in14 (1'b0),                                   // (terminated)
		.reset_in15     (1'b0),                                   // (terminated)
		.reset_req_in15 (1'b0)                                    // (terminated)
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS          (1),
		.OUTPUT_RESET_SYNC_EDGES   ("deassert"),
		.SYNC_DEPTH                (2),
		.RESET_REQUEST_PRESENT     (1),
		.RESET_REQ_WAIT_TIME       (1),
		.MIN_RST_ASSERTION_TIME    (3),
		.RESET_REQ_EARLY_DSRT_TIME (1),
		.USE_RESET_REQUEST_IN0     (0),
		.USE_RESET_REQUEST_IN1     (0),
		.USE_RESET_REQUEST_IN2     (0),
		.USE_RESET_REQUEST_IN3     (0),
		.USE_RESET_REQUEST_IN4     (0),
		.USE_RESET_REQUEST_IN5     (0),
		.USE_RESET_REQUEST_IN6     (0),
		.USE_RESET_REQUEST_IN7     (0),
		.USE_RESET_REQUEST_IN8     (0),
		.USE_RESET_REQUEST_IN9     (0),
		.USE_RESET_REQUEST_IN10    (0),
		.USE_RESET_REQUEST_IN11    (0),
		.USE_RESET_REQUEST_IN12    (0),
		.USE_RESET_REQUEST_IN13    (0),
		.USE_RESET_REQUEST_IN14    (0),
		.USE_RESET_REQUEST_IN15    (0),
		.ADAPT_RESET_REQUEST       (0)
	) rst_controller_002 (
		.reset_in0      (~reset_reset_n),                         // reset_in0.reset
		.clk            (clk_clk),                                //       clk.clk
		.reset_out      (rst_controller_002_reset_out_reset),     // reset_out.reset
		.reset_req      (rst_controller_002_reset_out_reset_req), //          .reset_req
		.reset_req_in0  (1'b0),                                   // (terminated)
		.reset_in1      (1'b0),                                   // (terminated)
		.reset_req_in1  (1'b0),                                   // (terminated)
		.reset_in2      (1'b0),                                   // (terminated)
		.reset_req_in2  (1'b0),                                   // (terminated)
		.reset_in3      (1'b0),                                   // (terminated)
		.reset_req_in3  (1'b0),                                   // (terminated)
		.reset_in4      (1'b0),                                   // (terminated)
		.reset_req_in4  (1'b0),                                   // (terminated)
		.reset_in5      (1'b0),                                   // (terminated)
		.reset_req_in5  (1'b0),                                   // (terminated)
		.reset_in6      (1'b0),                                   // (terminated)
		.reset_req_in6  (1'b0),                                   // (terminated)
		.reset_in7      (1'b0),                                   // (terminated)
		.reset_req_in7  (1'b0),                                   // (terminated)
		.reset_in8      (1'b0),                                   // (terminated)
		.reset_req_in8  (1'b0),                                   // (terminated)
		.reset_in9      (1'b0),                                   // (terminated)
		.reset_req_in9  (1'b0),                                   // (terminated)
		.reset_in10     (1'b0),                                   // (terminated)
		.reset_req_in10 (1'b0),                                   // (terminated)
		.reset_in11     (1'b0),                                   // (terminated)
		.reset_req_in11 (1'b0),                                   // (terminated)
		.reset_in12     (1'b0),                                   // (terminated)
		.reset_req_in12 (1'b0),                                   // (terminated)
		.reset_in13     (1'b0),                                   // (terminated)
		.reset_req_in13 (1'b0),                                   // (terminated)
		.reset_in14     (1'b0),                                   // (terminated)
		.reset_req_in14 (1'b0),                                   // (terminated)
		.reset_in15     (1'b0),                                   // (terminated)
		.reset_req_in15 (1'b0)                                    // (terminated)
	);

endmodule
